LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_arith.all;
USE IEEE.std_logic_unsigned.all;


ENTITY display IS
	PORT (
		entrada: IN STD_LOGIC_VECTOR(5 downto 0);

		display_unidade,
		display_dezena: OUT STD_LOGIC_VECTOR(6 downto 0)
	);
END display;

ARCHITECTURE behavior OF display IS

SIGNAL displays_buffer: STD_LOGIC_VECTOR (13 DOWNTO 0);

BEGIN
	WITH entrada SELECT
		displays_buffer <=
			"10000001000000" WHEN "000000", -- 0
			"10000001111001" WHEN "000001", -- 1
			"10000000100100" WHEN "000010", -- 2
			"10000000110000" WHEN "000011", -- 3
			"10000000011001" WHEN "000100", -- 4
			"10000000010010" WHEN "000101", -- 5
			"10000000000010" WHEN "000110", -- 6
			"10000001111000" WHEN "000111", -- 7
			"10000000000000" WHEN "001000", -- 8
			"10000000010000" WHEN "001001", -- 9
			"11110011000000" WHEN "001010", -- 10
			"11110011111001" WHEN "001011", -- 11
			"11110010100100" WHEN "001100", -- 12
			"11110010110000" WHEN "001101", -- 13
			"11110010011001" WHEN "001110", -- 14
			"11110010010010" WHEN "001111", -- 15
			"11110010000010" WHEN "010000", -- 16
			"11110011111000" WHEN "010001", -- 17
			"11110010000000" WHEN "010010", -- 18
			"11110010010000" WHEN "010011", -- 19
			"01001001000000" WHEN "010100", -- 20
			"01001001111001" WHEN "010101", -- 21
			"01001000100100" WHEN "010110", -- 22
			"01001000110000" WHEN "010111", -- 23
			"01001000011001" WHEN "011000", -- 24
			"01001000010010" WHEN "011001", -- 25
			"01001000000010" WHEN "011010", -- 26
			"01001001111000" WHEN "011011", -- 27
			"01001000000000" WHEN "011100", -- 28
			"01001000010000" WHEN "011101", -- 29
			"01100001000000" WHEN "011110", -- 30
			"01100001111001" WHEN "011111", -- 31
			"01100000100100" WHEN "100000", -- 32
			"01100000110000" WHEN "100001", -- 33
			"01100000011001" WHEN "100010", -- 34
			"01100000010010" WHEN "100011", -- 35
			"01100000000010" WHEN "100100", -- 36
			"01100001111000" WHEN "100101", -- 37
			"01100000000000" WHEN "100110", -- 38
			"01100000010000" WHEN "100111", -- 39
			"00110011000000" WHEN "101000", -- 40
			"00110011111001" WHEN "101001", -- 41
			"00110010100100" WHEN "101010", -- 42
			"00110010110000" WHEN "101011", -- 43
			"00110010011001" WHEN "101100", -- 44
			"00110010010010" WHEN "101101", -- 45
			"00110010000010" WHEN "101110", -- 46
			"00110011111000" WHEN "101111", -- 47
			"00110010000000" WHEN "110000", -- 48
			"00110010010000" WHEN "110001", -- 49
			"00100101000000" WHEN "110010", -- 50
			"00100101111001" WHEN "110011", -- 51
			"00100100100100" WHEN "110100", -- 52
			"00100100110000" WHEN "110101", -- 53
			"00100100011001" WHEN "110110", -- 54
			"00100100010010" WHEN "110111", -- 55
			"00100100000010" WHEN "111000", -- 56
			"00100101111000" WHEN "111001", -- 57
			"00100100000000" WHEN "111010", -- 58
			"00100100010000" WHEN "111011", -- 59
			"00000101000000" WHEN "111100", -- 60
			"00000101111001" WHEN "111101", -- 61
			"00000100100100" WHEN "111110", -- 62
			"00000100110000" WHEN "111111", -- 63
			"01111110111111" WHEN OTHERS;

	display_unidade <= displays_buffer(6 DOWNTO 0);
	display_dezena <= displays_buffer(13 DOWNTO 7);
END behavior;
